/home/runner/.cache/pip/pool/3a/ff/8b/d2ea50bc4cb88b8a1b64071929a20a49a72dccf5200e7aa54a9e3ee992